library verilog;
use verilog.vl_types.all;
entity testbench_fibonacci is
end testbench_fibonacci;
