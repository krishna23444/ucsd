// Platform Express Verilog testbench template
/**********************************************************************/
/*                    Px Generated File                               */
/*              Platform Express, Version 3.3.1 (BuildId: 200607071143)*/
/*              System Level Engineering Division                     */
/*              Mentor Graphics Corporation                           */
/*                                                                    */
/* Generated on: February 18, 2007 7:18:40 PM PST                     */
/* Generated by: saumya                                               */
/* Generated Top Level HDL                                            */
/**********************************************************************/



`timescale 1ns/1ps



// Testbench module
module pxdefault_tb;

// Signal Declaration
// 
// Signal Declaration for Component: test3_1
// 
    reg                  pxGen_ahb_1_HCLK;
    reg                  pxGen_ahb_1_HRESETn;
    reg                  pxGen_AHB_1_ambaAHB_HCLK;
    reg                  pxGen_AHB_1_ambaAHB_HRESETn;




// Component instantiation
// 
// Component: test3_1 Instantiation
// 

// 
//  Default value assignement for signals
// 
test3  test3_1(
    .test3_ahb_1_HCLK         (pxGen_ahb_1_HCLK),
    .test3_ahb_1_HRESETn      (pxGen_ahb_1_HRESETn),
    .test3_AHB_1_ambaAHB_HCLK (pxGen_AHB_1_ambaAHB_HCLK),
    .test3_AHB_1_ambaAHB_HRESETn(pxGen_AHB_1_ambaAHB_HRESETn) 
    );
// 
// Clock Driver ahb_1_HCLK

always begin
    pxGen_ahb_1_HCLK = 1'b1;
    #10.0 pxGen_ahb_1_HCLK = 1'b0;
    #20.0 pxGen_ahb_1_HCLK = 1'b1;
    #10.0 ;
end

// 
// Clock Driver AHB_1_ambaAHB_HCLK

always begin
    pxGen_AHB_1_ambaAHB_HCLK = 1'b1;
    #10.0 pxGen_AHB_1_ambaAHB_HCLK = 1'b0;
    #20.0 pxGen_AHB_1_ambaAHB_HCLK = 1'b1;
    #10.0 ;
end

// 
// Reset Drivers 

initial begin
    pxGen_ahb_1_HRESETn = 1'b1;
    #40.0 pxGen_ahb_1_HRESETn = 1'b0;
//    #24.0 pxGen_ahb_1_HRESETn = 1'b0;
    #800.0 pxGen_ahb_1_HRESETn = 1'b1;
end
initial begin
    pxGen_AHB_1_ambaAHB_HRESETn = 1'b1;
    #40.0 pxGen_AHB_1_ambaAHB_HRESETn = 1'b0;
//    #24.0 pxGen_AHB_1_ambaAHB_HRESETn = 1'b0;
    #800.0 pxGen_AHB_1_ambaAHB_HRESETn = 1'b1;
end




//
// VerificationIP instantiation
//
//@VerificationIP@

endmodule
